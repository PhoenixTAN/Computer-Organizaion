LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
ENTITY My16x8MUX IS
 PORT(
		--CLK: IN STD_LOGIC;
		Sout: IN STD_LOGIC;
		input: IN STD_LOGIC_VECTOR( 15 DOWNTO 0 );
		S: BUFFER STD_LOGIC_VECTOR( 7 DOWNTO 0 )
		);
END ENTITY My16x8MUX;

ARCHITECTURE TEST OF My16x8MUX IS
	SIGNAL Sel: STD_LOGIC;
BEGIN
	PROCESS(Sout)
	BEGIN
	--IF CLK'EVENT AND CLK = '1' THEN
		Sel <= Sout;
		IF SEL = '0' THEN			
			S <= input( 7 DOWNTO 0 );
		ELSIF Sout = '1' THEN
			S <= input( 15 DOWNTO 8 );
		END IF;
	--END IF;
	END PROCESS;
		
END ARCHITECTURE TEST;
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
ENTITY Adder_4 IS
	PORT(Ain,Bin,Cin: IN STD_LOGIC;
		Sum,Cout: out STD_LOGIC);
END Adder_4;

ARCHITECTURE rtl of Adder_4 IS	
	SIGNAL S: STD_LOGIC_VECTOR( 1 DOWNTO 0 );
BEGIN	
	S <= '0' & Ain + Bin + Cin;
	Sum <= S(0);
	Cout <= S(1);
END rtl;
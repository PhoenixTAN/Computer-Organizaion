LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
ENTITY My8x4MUX IS
 PORT(
		CLK: IN STD_LOGIC;
		Sout: IN STD_LOGIC;
		input: IN STD_LOGIC_VECTOR( 15 DOWNTO 0 );
		S: OUT STD_LOGIC_VECTOR( 7 DOWNTO 0 )
		);
END ENTITY My8x4MUX;

ARCHITECTURE TEST OF My8x4MUX IS
	SIGNAL Sel: STD_LOGIC;
BEGIN
	PROCESS(CLK)
	BEGIN
	IF CLK'EVENT AND CLK = '1' THEN
		Sel <= Sout;
		IF Sel = '0' THEN			
			S <= input( 7 DOWNTO 0 );
		ELSIF Sel = '1' THEN
			S <= input( 15 DOWNTO 8 );
		END IF;
	END IF;
	END PROCESS;
		
END ARCHITECTURE TEST;